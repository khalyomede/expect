module expect

pub struct Expectation[T] {
    actual_value T
}
